----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:38:22 09/12/2006 
-- Design Name: 
-- Module Name:    RAM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

library UNISIM;
use UNISIM.VComponents.all;

entity RAM is
  port (
    address : in  std_logic_vector (11 downto 0);
    clock   : in  std_logic;
    dataIn  : in  std_logic_vector (3 downto 0);
    dataOut : out std_logic_vector (3 downto 0);
    wrEn    : in  std_logic
    );

end RAM;

architecture Behavioral of RAM is

  signal SSR : std_logic;

begin

  -- RAMB16_S4: Virtex-II/II-Pro, Spartan-3/3E 4k x 4 Single-Port RAM
  -- Xilinx  HDL Language Template version 8.1i

  RAM_0 : RAMB16_S4
    generic map (
      INIT       => X"0",               --  Value of output RAM registers at startup
      SRVAL      => X"0",               --  Ouput value upon SSR assertion
      write_mode => "WRITE_FIRST",      --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      -- The following INIT_xx declarations specify the initial contents of the RAM
      -- Address 0 to 1023
      INIT_00    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F    => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 1024 to 2047
      INIT_10    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F    => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 2048 to 3071
      INIT_20    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F    => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 3072 to 4095
      INIT_30    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E    => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F    => X"0000000000000000000000000000000000000000000000000000000000000000")
    port map (
      DO         => dataOut,            -- 4-bit Data Output
      ADDR       => address,            -- 12-bit Address Input
      CLK        => clock,              -- Clock
      DI         => dataIn,             -- 4-bit Data Input
      EN         => '1',                -- RAM Enable Input
      SSR        => SSR,                -- Synchronous Set/Reset Input
      WE         => wrEn                -- Write Enable Input
      );

  -- End of RAMB16_S4_inst instantiation

end Behavioral;
